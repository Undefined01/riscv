`include "../common.v"

module mem(
);

	always @(*);

endmodule
